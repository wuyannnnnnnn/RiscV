module inst_fetch #(
    
)
(
    input   wire                     clk_i,
    input   wire                     rst_n_i,
);

always_ff @( posedge clk_i ) begin : blockName
    
end

endmodule
