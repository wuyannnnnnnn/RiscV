module core (
    input   wire                        clk_i,
    input   wire                        rst_n_i,

    
);
    
endmodule