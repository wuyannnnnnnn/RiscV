module id #(
    parameters
) (
    ports
);
    
endmodule